library ieee;
use ieee.std_logic_1164.all;

entity Controller is
    port (
        i_CLK : in std_logic;
        i_RST : in std_logic
    );
end entity;